module wallace(a,b,prod);
input [15:0] A;
input [15:0] B;
output[31:0] prod;
wire [15:0] p [15:0];
wire [20:0]s;
wire [20:0]c;
generate 
for(i=0;i<16;i++)
begin
assign p[i]= A & {16{B[i]}};
end
endgenerate

assign prod[0] = p[0][0];

generate 
for(i=0;i<16;i++)
begin
assign prod[i+1] = s[i];
end
endgenerate

ha ha1(p[0][1],p[1][0],s[0],c[0]);
fa fa1(p[0][2],p[1][1],p[2][0],s[1],c[1]);
fa fa2(p[0][3],p[1][2],p[2][1],s[2],c[2]);
fa fa3(p[0][4],p[1][3],p[2][2],s[3],c[3]);
fa fa4(p[0][5],p[1][4],p[2][3],s[4],c[4]);
fa fa5(p[0][6],p[1][5],p[2][4],s[5],c[5]);
fa fa6(p[0][7],p[1][6],p[2][5],s[6],c[6]);
fa fa7(p[0][8],p[1][7],p[2][6],s[7],c[7]);
fa fa8(p[0][9],p[1][8],p[2][7],s[8],c[8]);
fa fa9(p[0][10],p[1][9],p[2][8],s[9],c[9]);
fa fa10(p[0][11],p[1][10],p[2][9],s[10],c[10]);
fa fa11(p[0][12],p[1][11],p[2][10],s[11],c[11]);
fa fa12(p[0][13],p[1][12],p[2][11],s[12],c[12]);
fa fa13(p[0][14],p[1][13],p[2][12],s[13],c[13]);
fa fa14(p[0][15],p[1][14],p[2][13],s[14],c[14]);
fa fa15(p[1][15],p[2][14],p[3][13],s[15],c[15]);
fa fa16(p[2][15],p[3][14],p[4][13],s[16],c[16]);
fa fa17(p[3][15],p[4][14],p[5][13],s[17],c[17]);
fa fa18(p[4][15],p[5][14],p[6][13],s[18],c[18]);
fa fa19(p[5][15],p[6][14],p[7][13],s[19],c[19]);
fa fa20(p[6][15],p[7][14],p[8][13],s[20],c[20]);
fa fa21(p[7][15],p[8][14],p[9][13],s[21],c[21]);
fa fa22(p[8][15],p[9][14],p[10][13],s[22],c[22]);
fa fa23(p[9][15],p[10][14],p[11][13],s[23],c[23]);
fa fa24(p[10][15],p[11][14],p[12][13],s[24],c[24]);
fa fa25(p[11][15],p[12][14],p[13][13],s[25],c[25]);
fa fa26(p[12][15],p[13][14],p[14][13],s[26],c[26]);
fa fa27(p[13][15],p[14][14],p[15][13],s[27],c[27]);
ha ha28(p[14][15],p[15][14],s[28],c[28]);


ha ha30(c[0],s[1],s[29],c[29]);
fa fa31(p[3][0],c[1],s[2],s[30],c[30]);
fa fa31(p[3][1],c[2],s[3],s[31],c[31]);
fa fa32(p[3][2],c[3],s[4],s[32],c[32]);
fa fa33(p[3][3],c[4],s[5],s[33],c[33]);
fa fa34(p[3][4],c[5],s[6],s[34],c[34]);
fa fa35(p[3][5],c[6],s[7],s[35],c[35]);
fa fa36(p[3][6],c[7],s[8],s[36],c[36]);
fa fa37(p[3][7],c[8],s[9],s[37],c[37]);
fa fa38(p[3][8],c[9],s[10],s[38],c[38]);
fa fa39(p[3][9],c[10],s[11],s[39],c[39]);
fa fa40(p[3][10],c[11],s[12],s[40],c[40]);
fa fa41(p[3][11],c[12],s[13],s[41],c[41]);
fa fa42(p[3][12],c[13],s[14],s[42],c[42]);

fa fa43(p[4][12],c[14],s[15],s[43],c[43]);
fa fa44(p[5][12],c[15],s[16],s[44],c[44]);
fa fa45(p[6][12],c[16],s[17],s[45],c[45]);
fa fa46(p[7][12],c[17],s[18],s[46],c[46]);
fa fa47(p[8][12],c[18],s[19],s[47],c[47]);
fa fa48(p[9][12],c[19],s[20],s[48],c[48]);
fa fa49(p[10][12],c[20],s[21],s[49],c[49]);
fa fa50(p[11][12],c[21],s[22],s[50],c[50]);
fa fa51(p[12][12],c[22],s[23],s[51],c[51]);





fa fa52(p[13][13],c[23],s[24],s[52],c[52]);
fa fa53(p[12][13],c[22],s[23],s[51],c[51]);
fa fa54(p[11][13],c[21],s[22],s[50],c[50]);
fa fa55(p[12][13],c[22],s[23],s[51],c[51]);








