module shifter(in,shift,out);
input in[9:0],shift;
output out;


